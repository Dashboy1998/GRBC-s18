use work.word.all;

package DoubleQWord is 
	type DQWord is array (3 downto 0) of word;
end DoubleQWord;