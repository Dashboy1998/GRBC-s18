library ieee;
use ieee.std_logic_1164.all;

package byte is
	subtype byte is std_logic_vector(7 downto 0);				  
end byte;
