use work.byte.all;

package word is
	type word is array (0 to 3) of byte;
end word;