use work.byte.all;

package LUT2_array is
	type array_512 is array (0 to 511) of byte;
end LUT2_array;