use work.byte.all;

package LUT_array is
	type array_256 is array (0 to 255) of byte;
end LUT_array;